----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:43:47 04/08/2016 
-- Design Name: 
-- Module Name:    Division - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Division is
	generic(
		n : integer := 8;
		m : integer := 8
		);
	port(
		RST : in std_logic;
		CLK : in std_logic;
		A   
end Division;

architecture Behavioral of Division is

begin


end Behavioral;

